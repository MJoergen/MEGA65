library ieee;
use ieee.std_logic_1164.all;

package bitmap_pkg is
    type bitmap_t is array(0 to 255) of std_logic_vector(1 downto 0);

    constant bitmap_queen : bitmap_t := (
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","00","01","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","01","00","01","00","01","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","01","00","00","01","00","00","00","00",
        "00","00","00","00","00","00","01","00","01","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","00","01","00","01","00","01","00","00","00","00","00",
        "00","00","00","00","00","01","00","00","01","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","01","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","01","00","01","00","01","00","00","00","00",
        "00","00","00","00","00","00","01","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00");

    constant bitmap_grey : bitmap_t := (
        "01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
        "00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
        "01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
        "00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
        "01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
        "00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
        "01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
        "00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
        "01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
        "00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
        "01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
        "00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
        "01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
        "00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01",
        "01","00","01","00","01","00","01","00","01","00","01","00","01","00","01","00",
        "00","01","00","01","00","01","00","01","00","01","00","01","00","01","00","01");

    constant bitmap_0 : bitmap_t := (
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","00","01","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","00","01","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00");

    constant bitmap_1 : bitmap_t := (
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","01","01","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","01","01","01","01","01","01","01","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00");

    constant bitmap_2 : bitmap_t := (
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","00","01","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","01","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","01","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","01","01","01","01","01","01","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00");

    constant bitmap_3 : bitmap_t := (
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","01","01","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","01","01","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00");

    constant bitmap_4 : bitmap_t := (
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","01","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","01","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","01","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","01","01","01","01","01","01","01","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","01","01","01","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00");

    constant bitmap_5 : bitmap_t := (
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","01","01","01","01","01","01","00","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","01","01","01","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","01","01","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00");

    constant bitmap_6 : bitmap_t := (
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00",
        "00","00","00","00","00","00","00","01","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","01","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","01","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","01","00","01","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","01","01","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","00","01","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00");

    constant bitmap_7 : bitmap_t := (
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","01","01","01","01","01","01","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","01","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","01","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00");

    constant bitmap_8 : bitmap_t := (
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","00","01","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","00","01","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","00","01","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","00","01","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00");

    constant bitmap_9 : bitmap_t := (
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","00","01","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","00","01","00","00","00","01","01","00","00","00","00",
        "00","00","00","00","00","00","00","01","01","01","00","01","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00");

end package bitmap_pkg;

