library ieee;
   use ieee.std_logic_1164.all;

package bitmap_pkg is

   type     bitmap_type is array(0 to 255) of std_logic_vector(1 downto 0);

   constant C_BITMAP_0 : bitmap_type := (
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00");

   constant C_BITMAP_1 : bitmap_type := (
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "01", "00", "01", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00");

   constant C_BITMAP_2 : bitmap_type := (
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00");

   constant C_BITMAP_3 : bitmap_type := (
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00");

   constant C_BITMAP_4 : bitmap_type := (
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00");

   constant C_BITMAP_5 : bitmap_type := (
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "01", "01", "01", "01", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00");

   constant C_BITMAP_6 : bitmap_type := (
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00");

   constant C_BITMAP_7 : bitmap_type := (
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "01", "01", "01", "01", "01", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00");

   constant C_BITMAP_8 : bitmap_type := (
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00");

   constant C_BITMAP_9 : bitmap_type := (
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "01", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "01", "01", "01", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "01", "01", "01", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00",
                                           "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00");

end package bitmap_pkg;

